/*
DESCRIPTION

NOTES

TODO

*/

module example #(

)(

);

/**********
 * Internal Signals
**********/
/**********
 * Glue Logic 
 **********/
/**********
 * Synchronous Logic
 **********/
/**********
 * Glue Logic 
 **********/
/**********
 * Components
 **********/
/**********
 * Output Combinatorial Logic
 **********/
endmodule